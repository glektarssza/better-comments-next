-- ! comment
